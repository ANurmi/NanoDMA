module ndma_write_mgr #()();
endmodule : ndma_write_mgr
