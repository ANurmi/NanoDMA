module ndma_read_mgr #()();
endmodule : ndma_read_mgr
