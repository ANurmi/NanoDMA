module ndma #()();



endmodule : ndma
