module ndma_write_mgr #()(
  input  logic        clk_i,
  input  logic        rst_ni,
  input  logic [31:0] addr_i
);
endmodule : ndma_write_mgr
